
module mod1_top;
    mod1 mod1_inst();

    initial begin
        $display("Hello World!");
        $finish;
    end

endmodule
