
module mod1;

endmodule