
module err_syn;

abc;

endmddule

