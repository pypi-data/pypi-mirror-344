`include "uvm_macros.svh"

module top;

initial begin
    $display("Hello World!");
end

endmodule

