
module top;

    mod1 u_mod1();

    initial begin
        $display("Hello World!");
        $finish;
    end

endmodule